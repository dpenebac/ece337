// $Id: $
// File name:   tb_mealy.sv
// Created:     2/14/2022
// Author:      Dorien Penebacker
// Lab Section: 337-09
// Version:     1.0  Initial Design Entry
// Description: TestBench for Mealy Machine 1101 Detector
