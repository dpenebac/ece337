// $Id: $
// File name:   tb_adder_8bit.sv
// Created:     1/22/2022
// Author:      Dorien Penebacker
// Lab Section: 337-09
// Version:     1.0  Initial Design Entry
// Description: Test bench for adder_8bit
