// $Id: $
// File name:   adder_nbit.sv
// Created:     1/22/2022
// Author:      Dorien Penebacker
// Lab Section: 337-09
// Version:     1.0  Initial Design Entry
// Description: Parameterized Ripple Carry Adder
